-- Source: https://www.fpga4student.com/2018/08/basys-3-fpga-ov7670-camera.html
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity Address_Generator is
    Port ( 	CLK25,enable : in  STD_LOGIC;								-- horloge de 25 MHz et signal d'activation respectivement
            rst          : in STD_LOGIC;
            rez_160x120  : IN std_logic;
            rez_320x240  : IN std_logic;
            vsync        : in  STD_LOGIC;
				address 		 : out STD_LOGIC_VECTOR (18 downto 0));	-- adresse g�n�r�
end Address_Generator;

architecture Behavioral of Address_Generator is
   signal val: STD_LOGIC_VECTOR(address'range):= (others => '0');		-- signal intermidiaire
begin
	address <= val;																		-- adresse g�n�r�

	process(CLK25)
		begin
            if rising_edge(CLK25) then
                if rst = '1' then
                    val <= (others => '0');
                else
                    if (enable='1') then													-- si enable = 0 on arrete la g�n�ration d'adresses
                       if rez_160x120 = '1' then
                          if (val < 160*120) then										-- si l'espace m�moire est balay� compl�tement				
                             val <= val + 1 ;
                          end if;
                       elsif rez_320x240 = '1' then
                          if (val < 320*240) then										-- si l'espace m�moire est balay� compl�tement				
                             val <= val + 1 ;
                          end if;
                       else
                          if (val < 640*480) then										-- si l'espace m�moire est balay� compl�tement				
                             val <= val + 1 ;
                          end if;
                       end if;
                        end if;
                    if vsync = '0' then 
                       val <= (others => '0');
                    end if;
                end if;
            end if;	
		end process;
end Behavioral;

